//------------------------------------------------------------------------------
// Definitions and macros for RISCV agent
//------------------------------------------------------------------------------
// This file contains definitions and macros used by the RISCV agent.
//
// Author: Gustavo Santiago
// Date  : June 2025
//------------------------------------------------------------------------------

`ifndef RISCV_DEFINES
`define RISCV_DEFINES

  `define RISCV_WIDTH 4 
  `define NO_OF_TRANSACTIONS 10

  `define P_DATA_WIDTH 32
  `define P_ADDR_WIDTH 10
  `define P_REG_ADDR_WIDTH 5
  `define P_IMEM_ADDR_WIDTH 9
  `define P_DMEM_ADDR_WIDTH 8

`endif
