
module mux4to1 (
    input  logic [31:0] in0,
    input  logic [31:0] in1,
    input  logic [31:0] in2,
    input  logic [31:0] in3,
    input  logic [1:0]  sel,
    output logic [31:0] out
);
 
    always_comb begin
    out = in0;
        case (sel)
            2'b01: out = in1;
            2'b10: out = in2;
            2'b11: out = in3;
        endcase
    end
 
endmodule
